module S_ROM(cnt, S);
    input [5:0] cnt;
    output reg [4:0] S;

    always @(*)
        case(cnt)
            6'd0: S = 5'd7;
            6'd1: S = 5'd12;
            6'd2: S = 5'd17;
            6'd3: S = 5'd22;
            6'd4: S = 5'd7;
            6'd5: S = 5'd12;
            6'd6: S = 5'd17;
            6'd7: S = 5'd22;
            6'd8: S = 5'd7;
            6'd9: S = 5'd12;
            6'd10: S = 5'd17;
            6'd11: S = 5'd22;
            6'd12: S = 5'd7;
            6'd13: S = 5'd12;
            6'd14: S = 5'd17;
            6'd15: S = 5'd22;
            6'd16: S = 5'd5;
            6'd17: S = 5'd9;
            6'd18: S = 5'd14;
            6'd19: S = 5'd20;
            6'd20: S = 5'd5;
            6'd21: S = 5'd9;
            6'd22: S = 5'd14;
            6'd23: S = 5'd20;
            6'd24: S = 5'd5;
            6'd25: S = 5'd9;
            6'd26: S = 5'd14;
            6'd27: S = 5'd20;
            6'd28: S = 5'd5;
            6'd29: S = 5'd9;
            6'd30: S = 5'd14;
            6'd31: S = 5'd20;
            6'd32: S = 5'd4;
            6'd33: S = 5'd11;
            6'd34: S = 5'd16;
            6'd35: S = 5'd23;
            6'd36: S = 5'd4;
            6'd37: S = 5'd11;
            6'd38: S = 5'd16;
            6'd39: S = 5'd23;
            6'd40: S = 5'd4;
            6'd41: S = 5'd11;
            6'd42: S = 5'd16;
            6'd43: S = 5'd23;
            6'd44: S = 5'd4;
            6'd45: S = 5'd11;
            6'd46: S = 5'd16;
            6'd47: S = 5'd23;
            6'd48: S = 5'd6;
            6'd49: S = 5'd10;
            6'd50: S = 5'd15;
            6'd51: S = 5'd21;
            6'd52: S = 5'd6;
            6'd53: S = 5'd10;
            6'd54: S = 5'd15;
            6'd55: S = 5'd21;
            6'd56: S = 5'd6;
            6'd57: S = 5'd10;
            6'd58: S = 5'd15;
            6'd59: S = 5'd21;
            6'd60: S = 5'd6;
            6'd61: S = 5'd10;
            6'd62: S = 5'd15;
            6'd63: S = 5'd21;
        endcase
endmodule 
module hex15(x, y);
	input [3:0]x;
	output reg [6:0]y;
	
	always @(*) begin
		case(x) 
			4'b0000:y = 7'b1000000;
			4'b0001:y = 7'b1111001;
			4'b0010:y = 7'b0100100;
			4'b0011:y = 7'b0110000;
			4'b0100:y = 7'b0011001;
			4'b0101:y = 7'b0010010;
			4'b0110:y = 7'b0000010;
			4'b0111:y = 7'b1111000;
			4'b1000:y = 7'b0000000;
			4'b1001:y = 7'b0010000;
			4'b1010:y = 7'b0001000;
			4'b1011:y = 7'b0000011;
			4'b1100:y = 7'b1000110;
			4'b1101:y = 7'b0100001;
			4'b1110:y = 7'b0000110;
			4'b1111:y = 7'b0001110;
			default: y = 7'b1111111;
		endcase 
	end
	/*
		assign y[0] = (~x[3]&x[2]&~x[1]&~x[0])|(~x[3]&~x[2]&~x[1]&x[0])|(x[3]&x[2]&~x[1]&x[0])|(x[3]&~x[2]&x[1]&x[0]);
		assign y[1] = (~x[3]&x[2]&~x[1]&x[0])|(x[3]&x[2]&~x[0])|(x[3]&x[2]&x[1])|(x[2]&x[1]&~x[0])|(x[3]&x[1]&x[0]);
		assign y[2] = (~x[3]&~x[2]&x[1]&~x[0])|(x[3]&x[2]&~x[0])|(x[3]&x[2]&x[1]);
		assign y[3] = (~x[3]&~x[2]&~x[1]&x[0])|(x[2]&x[1]&x[0])|(x[3]&~x[2]&x[1]&~x[0])|(~x[3]&x[2]&~x[1]&~x[0]);
		assign y[4] = (~x[3]&x[2]&~x[1])|(~x[3]&x[0])|(x[3]&~x[2]&~x[1]&x[0]);
		assign y[5] = (~x[3]&~x[2]&(x[0]|x[1]))|(~x[3]&x[1]&x[0])|(x[3]&x[2]&~x[1]&x[0]);
		assign y[6] = (~x[3]&~x[2]&~x[1])|(x[3]&x[2]&~x[1]&~x[0])|(~x[3]&x[2]&x[1]&x[0]);
	*/
endmodule 
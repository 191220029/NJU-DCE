module string_commun();
input [7:0]ascii;
input [9:0] h_addr,
input [9:0] v_addr,
input read_clk, write_clk;
output [23:0]data;


endmodule;
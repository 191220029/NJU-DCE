module div_mod(h, v, map_h, map_v, mod9, mod16);
    input [9:0] h;
    input [9:0] v;

    output [4:0] map_v;
    output reg[6:0] map_h;
    output reg[3:0] mod9;
    output [3:0] mod16;

    //div9 div_nine(h, map_h, mod9);
    assign map_v = v[8:4];
    assign mod16 = v[3:0];
	 
	 always @*
    case(h)
        10'd0: begin map_h=7'd0; mod9=4'd0; end
        10'd1: begin map_h=7'd0; mod9=4'd1; end
        10'd2: begin map_h=7'd0; mod9=4'd2; end
        10'd3: begin map_h=7'd0; mod9=4'd3; end
        10'd4: begin map_h=7'd0; mod9=4'd4; end
        10'd5: begin map_h=7'd0; mod9=4'd5; end
        10'd6: begin map_h=7'd0; mod9=4'd6; end
        10'd7: begin map_h=7'd0; mod9=4'd7; end
        10'd8: begin map_h=7'd0; mod9=4'd8; end
        10'd9: begin map_h=7'd1; mod9=4'd0; end
        10'd10: begin map_h=7'd1; mod9=4'd1; end
        10'd11: begin map_h=7'd1; mod9=4'd2; end
        10'd12: begin map_h=7'd1; mod9=4'd3; end
        10'd13: begin map_h=7'd1; mod9=4'd4; end
        10'd14: begin map_h=7'd1; mod9=4'd5; end
        10'd15: begin map_h=7'd1; mod9=4'd6; end
        10'd16: begin map_h=7'd1; mod9=4'd7; end
        10'd17: begin map_h=7'd1; mod9=4'd8; end
        10'd18: begin map_h=7'd2; mod9=4'd0; end
        10'd19: begin map_h=7'd2; mod9=4'd1; end
        10'd20: begin map_h=7'd2; mod9=4'd2; end
        10'd21: begin map_h=7'd2; mod9=4'd3; end
        10'd22: begin map_h=7'd2; mod9=4'd4; end
        10'd23: begin map_h=7'd2; mod9=4'd5; end
        10'd24: begin map_h=7'd2; mod9=4'd6; end
        10'd25: begin map_h=7'd2; mod9=4'd7; end
        10'd26: begin map_h=7'd2; mod9=4'd8; end
        10'd27: begin map_h=7'd3; mod9=4'd0; end
        10'd28: begin map_h=7'd3; mod9=4'd1; end
        10'd29: begin map_h=7'd3; mod9=4'd2; end
        10'd30: begin map_h=7'd3; mod9=4'd3; end
        10'd31: begin map_h=7'd3; mod9=4'd4; end
        10'd32: begin map_h=7'd3; mod9=4'd5; end
        10'd33: begin map_h=7'd3; mod9=4'd6; end
        10'd34: begin map_h=7'd3; mod9=4'd7; end
        10'd35: begin map_h=7'd3; mod9=4'd8; end
        10'd36: begin map_h=7'd4; mod9=4'd0; end
        10'd37: begin map_h=7'd4; mod9=4'd1; end
        10'd38: begin map_h=7'd4; mod9=4'd2; end
        10'd39: begin map_h=7'd4; mod9=4'd3; end
        10'd40: begin map_h=7'd4; mod9=4'd4; end
        10'd41: begin map_h=7'd4; mod9=4'd5; end
        10'd42: begin map_h=7'd4; mod9=4'd6; end
        10'd43: begin map_h=7'd4; mod9=4'd7; end
        10'd44: begin map_h=7'd4; mod9=4'd8; end
        10'd45: begin map_h=7'd5; mod9=4'd0; end
        10'd46: begin map_h=7'd5; mod9=4'd1; end
        10'd47: begin map_h=7'd5; mod9=4'd2; end
        10'd48: begin map_h=7'd5; mod9=4'd3; end
        10'd49: begin map_h=7'd5; mod9=4'd4; end
        10'd50: begin map_h=7'd5; mod9=4'd5; end
        10'd51: begin map_h=7'd5; mod9=4'd6; end
        10'd52: begin map_h=7'd5; mod9=4'd7; end
        10'd53: begin map_h=7'd5; mod9=4'd8; end
        10'd54: begin map_h=7'd6; mod9=4'd0; end
        10'd55: begin map_h=7'd6; mod9=4'd1; end
        10'd56: begin map_h=7'd6; mod9=4'd2; end
        10'd57: begin map_h=7'd6; mod9=4'd3; end
        10'd58: begin map_h=7'd6; mod9=4'd4; end
        10'd59: begin map_h=7'd6; mod9=4'd5; end
        10'd60: begin map_h=7'd6; mod9=4'd6; end
        10'd61: begin map_h=7'd6; mod9=4'd7; end
        10'd62: begin map_h=7'd6; mod9=4'd8; end
        10'd63: begin map_h=7'd7; mod9=4'd0; end
        10'd64: begin map_h=7'd7; mod9=4'd1; end
        10'd65: begin map_h=7'd7; mod9=4'd2; end
        10'd66: begin map_h=7'd7; mod9=4'd3; end
        10'd67: begin map_h=7'd7; mod9=4'd4; end
        10'd68: begin map_h=7'd7; mod9=4'd5; end
        10'd69: begin map_h=7'd7; mod9=4'd6; end
        10'd70: begin map_h=7'd7; mod9=4'd7; end
        10'd71: begin map_h=7'd7; mod9=4'd8; end
        10'd72: begin map_h=7'd8; mod9=4'd0; end
        10'd73: begin map_h=7'd8; mod9=4'd1; end
        10'd74: begin map_h=7'd8; mod9=4'd2; end
        10'd75: begin map_h=7'd8; mod9=4'd3; end
        10'd76: begin map_h=7'd8; mod9=4'd4; end
        10'd77: begin map_h=7'd8; mod9=4'd5; end
        10'd78: begin map_h=7'd8; mod9=4'd6; end
        10'd79: begin map_h=7'd8; mod9=4'd7; end
        10'd80: begin map_h=7'd8; mod9=4'd8; end
        10'd81: begin map_h=7'd9; mod9=4'd0; end
        10'd82: begin map_h=7'd9; mod9=4'd1; end
        10'd83: begin map_h=7'd9; mod9=4'd2; end
        10'd84: begin map_h=7'd9; mod9=4'd3; end
        10'd85: begin map_h=7'd9; mod9=4'd4; end
        10'd86: begin map_h=7'd9; mod9=4'd5; end
        10'd87: begin map_h=7'd9; mod9=4'd6; end
        10'd88: begin map_h=7'd9; mod9=4'd7; end
        10'd89: begin map_h=7'd9; mod9=4'd8; end
        10'd90: begin map_h=7'd10; mod9=4'd0; end
        10'd91: begin map_h=7'd10; mod9=4'd1; end
        10'd92: begin map_h=7'd10; mod9=4'd2; end
        10'd93: begin map_h=7'd10; mod9=4'd3; end
        10'd94: begin map_h=7'd10; mod9=4'd4; end
        10'd95: begin map_h=7'd10; mod9=4'd5; end
        10'd96: begin map_h=7'd10; mod9=4'd6; end
        10'd97: begin map_h=7'd10; mod9=4'd7; end
        10'd98: begin map_h=7'd10; mod9=4'd8; end
        10'd99: begin map_h=7'd11; mod9=4'd0; end
        10'd100: begin map_h=7'd11; mod9=4'd1; end
        10'd101: begin map_h=7'd11; mod9=4'd2; end
        10'd102: begin map_h=7'd11; mod9=4'd3; end
        10'd103: begin map_h=7'd11; mod9=4'd4; end
        10'd104: begin map_h=7'd11; mod9=4'd5; end
        10'd105: begin map_h=7'd11; mod9=4'd6; end
        10'd106: begin map_h=7'd11; mod9=4'd7; end
        10'd107: begin map_h=7'd11; mod9=4'd8; end
        10'd108: begin map_h=7'd12; mod9=4'd0; end
        10'd109: begin map_h=7'd12; mod9=4'd1; end
        10'd110: begin map_h=7'd12; mod9=4'd2; end
        10'd111: begin map_h=7'd12; mod9=4'd3; end
        10'd112: begin map_h=7'd12; mod9=4'd4; end
        10'd113: begin map_h=7'd12; mod9=4'd5; end
        10'd114: begin map_h=7'd12; mod9=4'd6; end
        10'd115: begin map_h=7'd12; mod9=4'd7; end
        10'd116: begin map_h=7'd12; mod9=4'd8; end
        10'd117: begin map_h=7'd13; mod9=4'd0; end
        10'd118: begin map_h=7'd13; mod9=4'd1; end
        10'd119: begin map_h=7'd13; mod9=4'd2; end
        10'd120: begin map_h=7'd13; mod9=4'd3; end
        10'd121: begin map_h=7'd13; mod9=4'd4; end
        10'd122: begin map_h=7'd13; mod9=4'd5; end
        10'd123: begin map_h=7'd13; mod9=4'd6; end
        10'd124: begin map_h=7'd13; mod9=4'd7; end
        10'd125: begin map_h=7'd13; mod9=4'd8; end
        10'd126: begin map_h=7'd14; mod9=4'd0; end
        10'd127: begin map_h=7'd14; mod9=4'd1; end
        10'd128: begin map_h=7'd14; mod9=4'd2; end
        10'd129: begin map_h=7'd14; mod9=4'd3; end
        10'd130: begin map_h=7'd14; mod9=4'd4; end
        10'd131: begin map_h=7'd14; mod9=4'd5; end
        10'd132: begin map_h=7'd14; mod9=4'd6; end
        10'd133: begin map_h=7'd14; mod9=4'd7; end
        10'd134: begin map_h=7'd14; mod9=4'd8; end
        10'd135: begin map_h=7'd15; mod9=4'd0; end
        10'd136: begin map_h=7'd15; mod9=4'd1; end
        10'd137: begin map_h=7'd15; mod9=4'd2; end
        10'd138: begin map_h=7'd15; mod9=4'd3; end
        10'd139: begin map_h=7'd15; mod9=4'd4; end
        10'd140: begin map_h=7'd15; mod9=4'd5; end
        10'd141: begin map_h=7'd15; mod9=4'd6; end
        10'd142: begin map_h=7'd15; mod9=4'd7; end
        10'd143: begin map_h=7'd15; mod9=4'd8; end
        10'd144: begin map_h=7'd16; mod9=4'd0; end
        10'd145: begin map_h=7'd16; mod9=4'd1; end
        10'd146: begin map_h=7'd16; mod9=4'd2; end
        10'd147: begin map_h=7'd16; mod9=4'd3; end
        10'd148: begin map_h=7'd16; mod9=4'd4; end
        10'd149: begin map_h=7'd16; mod9=4'd5; end
        10'd150: begin map_h=7'd16; mod9=4'd6; end
        10'd151: begin map_h=7'd16; mod9=4'd7; end
        10'd152: begin map_h=7'd16; mod9=4'd8; end
        10'd153: begin map_h=7'd17; mod9=4'd0; end
        10'd154: begin map_h=7'd17; mod9=4'd1; end
        10'd155: begin map_h=7'd17; mod9=4'd2; end
        10'd156: begin map_h=7'd17; mod9=4'd3; end
        10'd157: begin map_h=7'd17; mod9=4'd4; end
        10'd158: begin map_h=7'd17; mod9=4'd5; end
        10'd159: begin map_h=7'd17; mod9=4'd6; end
        10'd160: begin map_h=7'd17; mod9=4'd7; end
        10'd161: begin map_h=7'd17; mod9=4'd8; end
        10'd162: begin map_h=7'd18; mod9=4'd0; end
        10'd163: begin map_h=7'd18; mod9=4'd1; end
        10'd164: begin map_h=7'd18; mod9=4'd2; end
        10'd165: begin map_h=7'd18; mod9=4'd3; end
        10'd166: begin map_h=7'd18; mod9=4'd4; end
        10'd167: begin map_h=7'd18; mod9=4'd5; end
        10'd168: begin map_h=7'd18; mod9=4'd6; end
        10'd169: begin map_h=7'd18; mod9=4'd7; end
        10'd170: begin map_h=7'd18; mod9=4'd8; end
        10'd171: begin map_h=7'd19; mod9=4'd0; end
        10'd172: begin map_h=7'd19; mod9=4'd1; end
        10'd173: begin map_h=7'd19; mod9=4'd2; end
        10'd174: begin map_h=7'd19; mod9=4'd3; end
        10'd175: begin map_h=7'd19; mod9=4'd4; end
        10'd176: begin map_h=7'd19; mod9=4'd5; end
        10'd177: begin map_h=7'd19; mod9=4'd6; end
        10'd178: begin map_h=7'd19; mod9=4'd7; end
        10'd179: begin map_h=7'd19; mod9=4'd8; end
        10'd180: begin map_h=7'd20; mod9=4'd0; end
        10'd181: begin map_h=7'd20; mod9=4'd1; end
        10'd182: begin map_h=7'd20; mod9=4'd2; end
        10'd183: begin map_h=7'd20; mod9=4'd3; end
        10'd184: begin map_h=7'd20; mod9=4'd4; end
        10'd185: begin map_h=7'd20; mod9=4'd5; end
        10'd186: begin map_h=7'd20; mod9=4'd6; end
        10'd187: begin map_h=7'd20; mod9=4'd7; end
        10'd188: begin map_h=7'd20; mod9=4'd8; end
        10'd189: begin map_h=7'd21; mod9=4'd0; end
        10'd190: begin map_h=7'd21; mod9=4'd1; end
        10'd191: begin map_h=7'd21; mod9=4'd2; end
        10'd192: begin map_h=7'd21; mod9=4'd3; end
        10'd193: begin map_h=7'd21; mod9=4'd4; end
        10'd194: begin map_h=7'd21; mod9=4'd5; end
        10'd195: begin map_h=7'd21; mod9=4'd6; end
        10'd196: begin map_h=7'd21; mod9=4'd7; end
        10'd197: begin map_h=7'd21; mod9=4'd8; end
        10'd198: begin map_h=7'd22; mod9=4'd0; end
        10'd199: begin map_h=7'd22; mod9=4'd1; end
        10'd200: begin map_h=7'd22; mod9=4'd2; end
        10'd201: begin map_h=7'd22; mod9=4'd3; end
        10'd202: begin map_h=7'd22; mod9=4'd4; end
        10'd203: begin map_h=7'd22; mod9=4'd5; end
        10'd204: begin map_h=7'd22; mod9=4'd6; end
        10'd205: begin map_h=7'd22; mod9=4'd7; end
        10'd206: begin map_h=7'd22; mod9=4'd8; end
        10'd207: begin map_h=7'd23; mod9=4'd0; end
        10'd208: begin map_h=7'd23; mod9=4'd1; end
        10'd209: begin map_h=7'd23; mod9=4'd2; end
        10'd210: begin map_h=7'd23; mod9=4'd3; end
        10'd211: begin map_h=7'd23; mod9=4'd4; end
        10'd212: begin map_h=7'd23; mod9=4'd5; end
        10'd213: begin map_h=7'd23; mod9=4'd6; end
        10'd214: begin map_h=7'd23; mod9=4'd7; end
        10'd215: begin map_h=7'd23; mod9=4'd8; end
        10'd216: begin map_h=7'd24; mod9=4'd0; end
        10'd217: begin map_h=7'd24; mod9=4'd1; end
        10'd218: begin map_h=7'd24; mod9=4'd2; end
        10'd219: begin map_h=7'd24; mod9=4'd3; end
        10'd220: begin map_h=7'd24; mod9=4'd4; end
        10'd221: begin map_h=7'd24; mod9=4'd5; end
        10'd222: begin map_h=7'd24; mod9=4'd6; end
        10'd223: begin map_h=7'd24; mod9=4'd7; end
        10'd224: begin map_h=7'd24; mod9=4'd8; end
        10'd225: begin map_h=7'd25; mod9=4'd0; end
        10'd226: begin map_h=7'd25; mod9=4'd1; end
        10'd227: begin map_h=7'd25; mod9=4'd2; end
        10'd228: begin map_h=7'd25; mod9=4'd3; end
        10'd229: begin map_h=7'd25; mod9=4'd4; end
        10'd230: begin map_h=7'd25; mod9=4'd5; end
        10'd231: begin map_h=7'd25; mod9=4'd6; end
        10'd232: begin map_h=7'd25; mod9=4'd7; end
        10'd233: begin map_h=7'd25; mod9=4'd8; end
        10'd234: begin map_h=7'd26; mod9=4'd0; end
        10'd235: begin map_h=7'd26; mod9=4'd1; end
        10'd236: begin map_h=7'd26; mod9=4'd2; end
        10'd237: begin map_h=7'd26; mod9=4'd3; end
        10'd238: begin map_h=7'd26; mod9=4'd4; end
        10'd239: begin map_h=7'd26; mod9=4'd5; end
        10'd240: begin map_h=7'd26; mod9=4'd6; end
        10'd241: begin map_h=7'd26; mod9=4'd7; end
        10'd242: begin map_h=7'd26; mod9=4'd8; end
        10'd243: begin map_h=7'd27; mod9=4'd0; end
        10'd244: begin map_h=7'd27; mod9=4'd1; end
        10'd245: begin map_h=7'd27; mod9=4'd2; end
        10'd246: begin map_h=7'd27; mod9=4'd3; end
        10'd247: begin map_h=7'd27; mod9=4'd4; end
        10'd248: begin map_h=7'd27; mod9=4'd5; end
        10'd249: begin map_h=7'd27; mod9=4'd6; end
        10'd250: begin map_h=7'd27; mod9=4'd7; end
        10'd251: begin map_h=7'd27; mod9=4'd8; end
        10'd252: begin map_h=7'd28; mod9=4'd0; end
        10'd253: begin map_h=7'd28; mod9=4'd1; end
        10'd254: begin map_h=7'd28; mod9=4'd2; end
        10'd255: begin map_h=7'd28; mod9=4'd3; end
        10'd256: begin map_h=7'd28; mod9=4'd4; end
        10'd257: begin map_h=7'd28; mod9=4'd5; end
        10'd258: begin map_h=7'd28; mod9=4'd6; end
        10'd259: begin map_h=7'd28; mod9=4'd7; end
        10'd260: begin map_h=7'd28; mod9=4'd8; end
        10'd261: begin map_h=7'd29; mod9=4'd0; end
        10'd262: begin map_h=7'd29; mod9=4'd1; end
        10'd263: begin map_h=7'd29; mod9=4'd2; end
        10'd264: begin map_h=7'd29; mod9=4'd3; end
        10'd265: begin map_h=7'd29; mod9=4'd4; end
        10'd266: begin map_h=7'd29; mod9=4'd5; end
        10'd267: begin map_h=7'd29; mod9=4'd6; end
        10'd268: begin map_h=7'd29; mod9=4'd7; end
        10'd269: begin map_h=7'd29; mod9=4'd8; end
        10'd270: begin map_h=7'd30; mod9=4'd0; end
        10'd271: begin map_h=7'd30; mod9=4'd1; end
        10'd272: begin map_h=7'd30; mod9=4'd2; end
        10'd273: begin map_h=7'd30; mod9=4'd3; end
        10'd274: begin map_h=7'd30; mod9=4'd4; end
        10'd275: begin map_h=7'd30; mod9=4'd5; end
        10'd276: begin map_h=7'd30; mod9=4'd6; end
        10'd277: begin map_h=7'd30; mod9=4'd7; end
        10'd278: begin map_h=7'd30; mod9=4'd8; end
        10'd279: begin map_h=7'd31; mod9=4'd0; end
        10'd280: begin map_h=7'd31; mod9=4'd1; end
        10'd281: begin map_h=7'd31; mod9=4'd2; end
        10'd282: begin map_h=7'd31; mod9=4'd3; end
        10'd283: begin map_h=7'd31; mod9=4'd4; end
        10'd284: begin map_h=7'd31; mod9=4'd5; end
        10'd285: begin map_h=7'd31; mod9=4'd6; end
        10'd286: begin map_h=7'd31; mod9=4'd7; end
        10'd287: begin map_h=7'd31; mod9=4'd8; end
        10'd288: begin map_h=7'd32; mod9=4'd0; end
        10'd289: begin map_h=7'd32; mod9=4'd1; end
        10'd290: begin map_h=7'd32; mod9=4'd2; end
        10'd291: begin map_h=7'd32; mod9=4'd3; end
        10'd292: begin map_h=7'd32; mod9=4'd4; end
        10'd293: begin map_h=7'd32; mod9=4'd5; end
        10'd294: begin map_h=7'd32; mod9=4'd6; end
        10'd295: begin map_h=7'd32; mod9=4'd7; end
        10'd296: begin map_h=7'd32; mod9=4'd8; end
        10'd297: begin map_h=7'd33; mod9=4'd0; end
        10'd298: begin map_h=7'd33; mod9=4'd1; end
        10'd299: begin map_h=7'd33; mod9=4'd2; end
        10'd300: begin map_h=7'd33; mod9=4'd3; end
        10'd301: begin map_h=7'd33; mod9=4'd4; end
        10'd302: begin map_h=7'd33; mod9=4'd5; end
        10'd303: begin map_h=7'd33; mod9=4'd6; end
        10'd304: begin map_h=7'd33; mod9=4'd7; end
        10'd305: begin map_h=7'd33; mod9=4'd8; end
        10'd306: begin map_h=7'd34; mod9=4'd0; end
        10'd307: begin map_h=7'd34; mod9=4'd1; end
        10'd308: begin map_h=7'd34; mod9=4'd2; end
        10'd309: begin map_h=7'd34; mod9=4'd3; end
        10'd310: begin map_h=7'd34; mod9=4'd4; end
        10'd311: begin map_h=7'd34; mod9=4'd5; end
        10'd312: begin map_h=7'd34; mod9=4'd6; end
        10'd313: begin map_h=7'd34; mod9=4'd7; end
        10'd314: begin map_h=7'd34; mod9=4'd8; end
        10'd315: begin map_h=7'd35; mod9=4'd0; end
        10'd316: begin map_h=7'd35; mod9=4'd1; end
        10'd317: begin map_h=7'd35; mod9=4'd2; end
        10'd318: begin map_h=7'd35; mod9=4'd3; end
        10'd319: begin map_h=7'd35; mod9=4'd4; end
        10'd320: begin map_h=7'd35; mod9=4'd5; end
        10'd321: begin map_h=7'd35; mod9=4'd6; end
        10'd322: begin map_h=7'd35; mod9=4'd7; end
        10'd323: begin map_h=7'd35; mod9=4'd8; end
        10'd324: begin map_h=7'd36; mod9=4'd0; end
        10'd325: begin map_h=7'd36; mod9=4'd1; end
        10'd326: begin map_h=7'd36; mod9=4'd2; end
        10'd327: begin map_h=7'd36; mod9=4'd3; end
        10'd328: begin map_h=7'd36; mod9=4'd4; end
        10'd329: begin map_h=7'd36; mod9=4'd5; end
        10'd330: begin map_h=7'd36; mod9=4'd6; end
        10'd331: begin map_h=7'd36; mod9=4'd7; end
        10'd332: begin map_h=7'd36; mod9=4'd8; end
        10'd333: begin map_h=7'd37; mod9=4'd0; end
        10'd334: begin map_h=7'd37; mod9=4'd1; end
        10'd335: begin map_h=7'd37; mod9=4'd2; end
        10'd336: begin map_h=7'd37; mod9=4'd3; end
        10'd337: begin map_h=7'd37; mod9=4'd4; end
        10'd338: begin map_h=7'd37; mod9=4'd5; end
        10'd339: begin map_h=7'd37; mod9=4'd6; end
        10'd340: begin map_h=7'd37; mod9=4'd7; end
        10'd341: begin map_h=7'd37; mod9=4'd8; end
        10'd342: begin map_h=7'd38; mod9=4'd0; end
        10'd343: begin map_h=7'd38; mod9=4'd1; end
        10'd344: begin map_h=7'd38; mod9=4'd2; end
        10'd345: begin map_h=7'd38; mod9=4'd3; end
        10'd346: begin map_h=7'd38; mod9=4'd4; end
        10'd347: begin map_h=7'd38; mod9=4'd5; end
        10'd348: begin map_h=7'd38; mod9=4'd6; end
        10'd349: begin map_h=7'd38; mod9=4'd7; end
        10'd350: begin map_h=7'd38; mod9=4'd8; end
        10'd351: begin map_h=7'd39; mod9=4'd0; end
        10'd352: begin map_h=7'd39; mod9=4'd1; end
        10'd353: begin map_h=7'd39; mod9=4'd2; end
        10'd354: begin map_h=7'd39; mod9=4'd3; end
        10'd355: begin map_h=7'd39; mod9=4'd4; end
        10'd356: begin map_h=7'd39; mod9=4'd5; end
        10'd357: begin map_h=7'd39; mod9=4'd6; end
        10'd358: begin map_h=7'd39; mod9=4'd7; end
        10'd359: begin map_h=7'd39; mod9=4'd8; end
        10'd360: begin map_h=7'd40; mod9=4'd0; end
        10'd361: begin map_h=7'd40; mod9=4'd1; end
        10'd362: begin map_h=7'd40; mod9=4'd2; end
        10'd363: begin map_h=7'd40; mod9=4'd3; end
        10'd364: begin map_h=7'd40; mod9=4'd4; end
        10'd365: begin map_h=7'd40; mod9=4'd5; end
        10'd366: begin map_h=7'd40; mod9=4'd6; end
        10'd367: begin map_h=7'd40; mod9=4'd7; end
        10'd368: begin map_h=7'd40; mod9=4'd8; end
        10'd369: begin map_h=7'd41; mod9=4'd0; end
        10'd370: begin map_h=7'd41; mod9=4'd1; end
        10'd371: begin map_h=7'd41; mod9=4'd2; end
        10'd372: begin map_h=7'd41; mod9=4'd3; end
        10'd373: begin map_h=7'd41; mod9=4'd4; end
        10'd374: begin map_h=7'd41; mod9=4'd5; end
        10'd375: begin map_h=7'd41; mod9=4'd6; end
        10'd376: begin map_h=7'd41; mod9=4'd7; end
        10'd377: begin map_h=7'd41; mod9=4'd8; end
        10'd378: begin map_h=7'd42; mod9=4'd0; end
        10'd379: begin map_h=7'd42; mod9=4'd1; end
        10'd380: begin map_h=7'd42; mod9=4'd2; end
        10'd381: begin map_h=7'd42; mod9=4'd3; end
        10'd382: begin map_h=7'd42; mod9=4'd4; end
        10'd383: begin map_h=7'd42; mod9=4'd5; end
        10'd384: begin map_h=7'd42; mod9=4'd6; end
        10'd385: begin map_h=7'd42; mod9=4'd7; end
        10'd386: begin map_h=7'd42; mod9=4'd8; end
        10'd387: begin map_h=7'd43; mod9=4'd0; end
        10'd388: begin map_h=7'd43; mod9=4'd1; end
        10'd389: begin map_h=7'd43; mod9=4'd2; end
        10'd390: begin map_h=7'd43; mod9=4'd3; end
        10'd391: begin map_h=7'd43; mod9=4'd4; end
        10'd392: begin map_h=7'd43; mod9=4'd5; end
        10'd393: begin map_h=7'd43; mod9=4'd6; end
        10'd394: begin map_h=7'd43; mod9=4'd7; end
        10'd395: begin map_h=7'd43; mod9=4'd8; end
        10'd396: begin map_h=7'd44; mod9=4'd0; end
        10'd397: begin map_h=7'd44; mod9=4'd1; end
        10'd398: begin map_h=7'd44; mod9=4'd2; end
        10'd399: begin map_h=7'd44; mod9=4'd3; end
        10'd400: begin map_h=7'd44; mod9=4'd4; end
        10'd401: begin map_h=7'd44; mod9=4'd5; end
        10'd402: begin map_h=7'd44; mod9=4'd6; end
        10'd403: begin map_h=7'd44; mod9=4'd7; end
        10'd404: begin map_h=7'd44; mod9=4'd8; end
        10'd405: begin map_h=7'd45; mod9=4'd0; end
        10'd406: begin map_h=7'd45; mod9=4'd1; end
        10'd407: begin map_h=7'd45; mod9=4'd2; end
        10'd408: begin map_h=7'd45; mod9=4'd3; end
        10'd409: begin map_h=7'd45; mod9=4'd4; end
        10'd410: begin map_h=7'd45; mod9=4'd5; end
        10'd411: begin map_h=7'd45; mod9=4'd6; end
        10'd412: begin map_h=7'd45; mod9=4'd7; end
        10'd413: begin map_h=7'd45; mod9=4'd8; end
        10'd414: begin map_h=7'd46; mod9=4'd0; end
        10'd415: begin map_h=7'd46; mod9=4'd1; end
        10'd416: begin map_h=7'd46; mod9=4'd2; end
        10'd417: begin map_h=7'd46; mod9=4'd3; end
        10'd418: begin map_h=7'd46; mod9=4'd4; end
        10'd419: begin map_h=7'd46; mod9=4'd5; end
        10'd420: begin map_h=7'd46; mod9=4'd6; end
        10'd421: begin map_h=7'd46; mod9=4'd7; end
        10'd422: begin map_h=7'd46; mod9=4'd8; end
        10'd423: begin map_h=7'd47; mod9=4'd0; end
        10'd424: begin map_h=7'd47; mod9=4'd1; end
        10'd425: begin map_h=7'd47; mod9=4'd2; end
        10'd426: begin map_h=7'd47; mod9=4'd3; end
        10'd427: begin map_h=7'd47; mod9=4'd4; end
        10'd428: begin map_h=7'd47; mod9=4'd5; end
        10'd429: begin map_h=7'd47; mod9=4'd6; end
        10'd430: begin map_h=7'd47; mod9=4'd7; end
        10'd431: begin map_h=7'd47; mod9=4'd8; end
        10'd432: begin map_h=7'd48; mod9=4'd0; end
        10'd433: begin map_h=7'd48; mod9=4'd1; end
        10'd434: begin map_h=7'd48; mod9=4'd2; end
        10'd435: begin map_h=7'd48; mod9=4'd3; end
        10'd436: begin map_h=7'd48; mod9=4'd4; end
        10'd437: begin map_h=7'd48; mod9=4'd5; end
        10'd438: begin map_h=7'd48; mod9=4'd6; end
        10'd439: begin map_h=7'd48; mod9=4'd7; end
        10'd440: begin map_h=7'd48; mod9=4'd8; end
        10'd441: begin map_h=7'd49; mod9=4'd0; end
        10'd442: begin map_h=7'd49; mod9=4'd1; end
        10'd443: begin map_h=7'd49; mod9=4'd2; end
        10'd444: begin map_h=7'd49; mod9=4'd3; end
        10'd445: begin map_h=7'd49; mod9=4'd4; end
        10'd446: begin map_h=7'd49; mod9=4'd5; end
        10'd447: begin map_h=7'd49; mod9=4'd6; end
        10'd448: begin map_h=7'd49; mod9=4'd7; end
        10'd449: begin map_h=7'd49; mod9=4'd8; end
        10'd450: begin map_h=7'd50; mod9=4'd0; end
        10'd451: begin map_h=7'd50; mod9=4'd1; end
        10'd452: begin map_h=7'd50; mod9=4'd2; end
        10'd453: begin map_h=7'd50; mod9=4'd3; end
        10'd454: begin map_h=7'd50; mod9=4'd4; end
        10'd455: begin map_h=7'd50; mod9=4'd5; end
        10'd456: begin map_h=7'd50; mod9=4'd6; end
        10'd457: begin map_h=7'd50; mod9=4'd7; end
        10'd458: begin map_h=7'd50; mod9=4'd8; end
        10'd459: begin map_h=7'd51; mod9=4'd0; end
        10'd460: begin map_h=7'd51; mod9=4'd1; end
        10'd461: begin map_h=7'd51; mod9=4'd2; end
        10'd462: begin map_h=7'd51; mod9=4'd3; end
        10'd463: begin map_h=7'd51; mod9=4'd4; end
        10'd464: begin map_h=7'd51; mod9=4'd5; end
        10'd465: begin map_h=7'd51; mod9=4'd6; end
        10'd466: begin map_h=7'd51; mod9=4'd7; end
        10'd467: begin map_h=7'd51; mod9=4'd8; end
        10'd468: begin map_h=7'd52; mod9=4'd0; end
        10'd469: begin map_h=7'd52; mod9=4'd1; end
        10'd470: begin map_h=7'd52; mod9=4'd2; end
        10'd471: begin map_h=7'd52; mod9=4'd3; end
        10'd472: begin map_h=7'd52; mod9=4'd4; end
        10'd473: begin map_h=7'd52; mod9=4'd5; end
        10'd474: begin map_h=7'd52; mod9=4'd6; end
        10'd475: begin map_h=7'd52; mod9=4'd7; end
        10'd476: begin map_h=7'd52; mod9=4'd8; end
        10'd477: begin map_h=7'd53; mod9=4'd0; end
        10'd478: begin map_h=7'd53; mod9=4'd1; end
        10'd479: begin map_h=7'd53; mod9=4'd2; end
        10'd480: begin map_h=7'd53; mod9=4'd3; end
        10'd481: begin map_h=7'd53; mod9=4'd4; end
        10'd482: begin map_h=7'd53; mod9=4'd5; end
        10'd483: begin map_h=7'd53; mod9=4'd6; end
        10'd484: begin map_h=7'd53; mod9=4'd7; end
        10'd485: begin map_h=7'd53; mod9=4'd8; end
        10'd486: begin map_h=7'd54; mod9=4'd0; end
        10'd487: begin map_h=7'd54; mod9=4'd1; end
        10'd488: begin map_h=7'd54; mod9=4'd2; end
        10'd489: begin map_h=7'd54; mod9=4'd3; end
        10'd490: begin map_h=7'd54; mod9=4'd4; end
        10'd491: begin map_h=7'd54; mod9=4'd5; end
        10'd492: begin map_h=7'd54; mod9=4'd6; end
        10'd493: begin map_h=7'd54; mod9=4'd7; end
        10'd494: begin map_h=7'd54; mod9=4'd8; end
        10'd495: begin map_h=7'd55; mod9=4'd0; end
        10'd496: begin map_h=7'd55; mod9=4'd1; end
        10'd497: begin map_h=7'd55; mod9=4'd2; end
        10'd498: begin map_h=7'd55; mod9=4'd3; end
        10'd499: begin map_h=7'd55; mod9=4'd4; end
        10'd500: begin map_h=7'd55; mod9=4'd5; end
        10'd501: begin map_h=7'd55; mod9=4'd6; end
        10'd502: begin map_h=7'd55; mod9=4'd7; end
        10'd503: begin map_h=7'd55; mod9=4'd8; end
        10'd504: begin map_h=7'd56; mod9=4'd0; end
        10'd505: begin map_h=7'd56; mod9=4'd1; end
        10'd506: begin map_h=7'd56; mod9=4'd2; end
        10'd507: begin map_h=7'd56; mod9=4'd3; end
        10'd508: begin map_h=7'd56; mod9=4'd4; end
        10'd509: begin map_h=7'd56; mod9=4'd5; end
        10'd510: begin map_h=7'd56; mod9=4'd6; end
        10'd511: begin map_h=7'd56; mod9=4'd7; end
        10'd512: begin map_h=7'd56; mod9=4'd8; end
        10'd513: begin map_h=7'd57; mod9=4'd0; end
        10'd514: begin map_h=7'd57; mod9=4'd1; end
        10'd515: begin map_h=7'd57; mod9=4'd2; end
        10'd516: begin map_h=7'd57; mod9=4'd3; end
        10'd517: begin map_h=7'd57; mod9=4'd4; end
        10'd518: begin map_h=7'd57; mod9=4'd5; end
        10'd519: begin map_h=7'd57; mod9=4'd6; end
        10'd520: begin map_h=7'd57; mod9=4'd7; end
        10'd521: begin map_h=7'd57; mod9=4'd8; end
        10'd522: begin map_h=7'd58; mod9=4'd0; end
        10'd523: begin map_h=7'd58; mod9=4'd1; end
        10'd524: begin map_h=7'd58; mod9=4'd2; end
        10'd525: begin map_h=7'd58; mod9=4'd3; end
        10'd526: begin map_h=7'd58; mod9=4'd4; end
        10'd527: begin map_h=7'd58; mod9=4'd5; end
        10'd528: begin map_h=7'd58; mod9=4'd6; end
        10'd529: begin map_h=7'd58; mod9=4'd7; end
        10'd530: begin map_h=7'd58; mod9=4'd8; end
        10'd531: begin map_h=7'd59; mod9=4'd0; end
        10'd532: begin map_h=7'd59; mod9=4'd1; end
        10'd533: begin map_h=7'd59; mod9=4'd2; end
        10'd534: begin map_h=7'd59; mod9=4'd3; end
        10'd535: begin map_h=7'd59; mod9=4'd4; end
        10'd536: begin map_h=7'd59; mod9=4'd5; end
        10'd537: begin map_h=7'd59; mod9=4'd6; end
        10'd538: begin map_h=7'd59; mod9=4'd7; end
        10'd539: begin map_h=7'd59; mod9=4'd8; end
        10'd540: begin map_h=7'd60; mod9=4'd0; end
        10'd541: begin map_h=7'd60; mod9=4'd1; end
        10'd542: begin map_h=7'd60; mod9=4'd2; end
        10'd543: begin map_h=7'd60; mod9=4'd3; end
        10'd544: begin map_h=7'd60; mod9=4'd4; end
        10'd545: begin map_h=7'd60; mod9=4'd5; end
        10'd546: begin map_h=7'd60; mod9=4'd6; end
        10'd547: begin map_h=7'd60; mod9=4'd7; end
        10'd548: begin map_h=7'd60; mod9=4'd8; end
        10'd549: begin map_h=7'd61; mod9=4'd0; end
        10'd550: begin map_h=7'd61; mod9=4'd1; end
        10'd551: begin map_h=7'd61; mod9=4'd2; end
        10'd552: begin map_h=7'd61; mod9=4'd3; end
        10'd553: begin map_h=7'd61; mod9=4'd4; end
        10'd554: begin map_h=7'd61; mod9=4'd5; end
        10'd555: begin map_h=7'd61; mod9=4'd6; end
        10'd556: begin map_h=7'd61; mod9=4'd7; end
        10'd557: begin map_h=7'd61; mod9=4'd8; end
        10'd558: begin map_h=7'd62; mod9=4'd0; end
        10'd559: begin map_h=7'd62; mod9=4'd1; end
        10'd560: begin map_h=7'd62; mod9=4'd2; end
        10'd561: begin map_h=7'd62; mod9=4'd3; end
        10'd562: begin map_h=7'd62; mod9=4'd4; end
        10'd563: begin map_h=7'd62; mod9=4'd5; end
        10'd564: begin map_h=7'd62; mod9=4'd6; end
        10'd565: begin map_h=7'd62; mod9=4'd7; end
        10'd566: begin map_h=7'd62; mod9=4'd8; end
        10'd567: begin map_h=7'd63; mod9=4'd0; end
        10'd568: begin map_h=7'd63; mod9=4'd1; end
        10'd569: begin map_h=7'd63; mod9=4'd2; end
        10'd570: begin map_h=7'd63; mod9=4'd3; end
        10'd571: begin map_h=7'd63; mod9=4'd4; end
        10'd572: begin map_h=7'd63; mod9=4'd5; end
        10'd573: begin map_h=7'd63; mod9=4'd6; end
        10'd574: begin map_h=7'd63; mod9=4'd7; end
        10'd575: begin map_h=7'd63; mod9=4'd8; end
        10'd576: begin map_h=7'd64; mod9=4'd0; end
        10'd577: begin map_h=7'd64; mod9=4'd1; end
        10'd578: begin map_h=7'd64; mod9=4'd2; end
        10'd579: begin map_h=7'd64; mod9=4'd3; end
        10'd580: begin map_h=7'd64; mod9=4'd4; end
        10'd581: begin map_h=7'd64; mod9=4'd5; end
        10'd582: begin map_h=7'd64; mod9=4'd6; end
        10'd583: begin map_h=7'd64; mod9=4'd7; end
        10'd584: begin map_h=7'd64; mod9=4'd8; end
        10'd585: begin map_h=7'd65; mod9=4'd0; end
        10'd586: begin map_h=7'd65; mod9=4'd1; end
        10'd587: begin map_h=7'd65; mod9=4'd2; end
        10'd588: begin map_h=7'd65; mod9=4'd3; end
        10'd589: begin map_h=7'd65; mod9=4'd4; end
        10'd590: begin map_h=7'd65; mod9=4'd5; end
        10'd591: begin map_h=7'd65; mod9=4'd6; end
        10'd592: begin map_h=7'd65; mod9=4'd7; end
        10'd593: begin map_h=7'd65; mod9=4'd8; end
        10'd594: begin map_h=7'd66; mod9=4'd0; end
        10'd595: begin map_h=7'd66; mod9=4'd1; end
        10'd596: begin map_h=7'd66; mod9=4'd2; end
        10'd597: begin map_h=7'd66; mod9=4'd3; end
        10'd598: begin map_h=7'd66; mod9=4'd4; end
        10'd599: begin map_h=7'd66; mod9=4'd5; end
        10'd600: begin map_h=7'd66; mod9=4'd6; end
        10'd601: begin map_h=7'd66; mod9=4'd7; end
        10'd602: begin map_h=7'd66; mod9=4'd8; end
        10'd603: begin map_h=7'd67; mod9=4'd0; end
        10'd604: begin map_h=7'd67; mod9=4'd1; end
        10'd605: begin map_h=7'd67; mod9=4'd2; end
        10'd606: begin map_h=7'd67; mod9=4'd3; end
        10'd607: begin map_h=7'd67; mod9=4'd4; end
        10'd608: begin map_h=7'd67; mod9=4'd5; end
        10'd609: begin map_h=7'd67; mod9=4'd6; end
        10'd610: begin map_h=7'd67; mod9=4'd7; end
        10'd611: begin map_h=7'd67; mod9=4'd8; end
        10'd612: begin map_h=7'd68; mod9=4'd0; end
        10'd613: begin map_h=7'd68; mod9=4'd1; end
        10'd614: begin map_h=7'd68; mod9=4'd2; end
        10'd615: begin map_h=7'd68; mod9=4'd3; end
        10'd616: begin map_h=7'd68; mod9=4'd4; end
        10'd617: begin map_h=7'd68; mod9=4'd5; end
        10'd618: begin map_h=7'd68; mod9=4'd6; end
        10'd619: begin map_h=7'd68; mod9=4'd7; end
        10'd620: begin map_h=7'd68; mod9=4'd8; end
        10'd621: begin map_h=7'd69; mod9=4'd0; end
        10'd622: begin map_h=7'd69; mod9=4'd1; end
        10'd623: begin map_h=7'd69; mod9=4'd2; end
        10'd624: begin map_h=7'd69; mod9=4'd3; end
        10'd625: begin map_h=7'd69; mod9=4'd4; end
        10'd626: begin map_h=7'd69; mod9=4'd5; end
        10'd627: begin map_h=7'd69; mod9=4'd6; end
        10'd628: begin map_h=7'd69; mod9=4'd7; end
        10'd629: begin map_h=7'd69; mod9=4'd8; end
        10'd630: begin map_h=7'd70; mod9=4'd0; end
        10'd631: begin map_h=7'd70; mod9=4'd1; end
        10'd632: begin map_h=7'd70; mod9=4'd2; end
        10'd633: begin map_h=7'd70; mod9=4'd3; end
        10'd634: begin map_h=7'd70; mod9=4'd4; end
        10'd635: begin map_h=7'd70; mod9=4'd5; end
        10'd636: begin map_h=7'd70; mod9=4'd6; end
        10'd637: begin map_h=7'd70; mod9=4'd7; end
        10'd638: begin map_h=7'd70; mod9=4'd8; end
        10'd639: begin map_h=7'd71; mod9=4'd0; end
        10'd640: begin map_h=7'd71; mod9=4'd1; end
        10'd641: begin map_h=7'd71; mod9=4'd2; end
        10'd642: begin map_h=7'd71; mod9=4'd3; end
        10'd643: begin map_h=7'd71; mod9=4'd4; end
        10'd644: begin map_h=7'd71; mod9=4'd5; end
        10'd645: begin map_h=7'd71; mod9=4'd6; end
        10'd646: begin map_h=7'd71; mod9=4'd7; end
        10'd647: begin map_h=7'd71; mod9=4'd8; end
        default: begin map_h = 7'd0; mod9 = 4'd0; end
    endcase
	 
endmodule

    